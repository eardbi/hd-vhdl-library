------------------------------------------------------------------------------
-- Title      : HDC Enhanced Package
-- Project    : Semester Thesis I
-------------------------------------------------------------------------------
-- File       : hdc_enhanced_pkg.vhd
-- Author     : Manuel Schmuck <schmucma@student.ethz.ch>
-- Company    : Integrated Systems Laboratory, ETH Zurich
-- Created    : 2017-09-30
-- Last update: 2018-01-02
-- Platform   : ModelSim (simulation), Vivado (synthesis)
-------------------------------------------------------------------------------
-- Description: Provides seed vectors and connectivity matrices for the
--              enhanced architecture.
-------------------------------------------------------------------------------
-- Copyright (c) 2017 Integrated Systems Laboratory, ETH Zurich
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author    Description
-- 2018        1.0      schmucma  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.hdc_pkg.all;

-------------------------------------------------------------------------------

package hdc_enhanced_pkg is

  -----------------------------------------------------------------------------
  -- Function Declarations
  -----------------------------------------------------------------------------
  

  -----------------------------------------------------------------------------
  -- Constant Declarations
  -----------------------------------------------------------------------------
  constant NHOT_LUT : std_logic_vector_array(0 to INPUT_QUANTIZATION-1)(0 to INPUT_QUANTIZATION-2) := (
		"00000000000000000000",
		"10000000000000000000",
		"11000000000000000000",
		"11100000000000000000",
		"11110000000000000000",
		"11111000000000000000",
		"11111100000000000000",
		"11111110000000000000",
		"11111111000000000000",
		"11111111100000000000",
		"11111111110000000000",
		"11111111111000000000",
		"11111111111100000000",
		"11111111111110000000",
		"11111111111111000000",
		"11111111111111100000",
		"11111111111111110000",
		"11111111111111111000",
		"11111111111111111100",
		"11111111111111111110",
		"11111111111111111111"
    );

  constant IM_SEED : hypervector(0 to HV_DIMENSION-1) := (
		"1001101110010101000100000101101111110110111101011000110110100011101010100100100100001011000110110110010101100001111100000110111111100101000000000010111011011110111010001011010011100100001001010011101011010011010110011101000001011111000001001101110100101111110101000111010000010110101110100110111000110000000001110010001110010100100010100111111001011011000000000000000000000100101110011000110101110100000010100111001110011111001100100100000100101001100101010110101010110101011000110110000100111001110001111011010001101100000100011111110000000111001111111110110111010011011101110101110100000000010100010010000101111011110111000110101100011110000011101101010111001111101010111101101110010010010100100011001000001010010101010001000001111010111010100111010110100011000101010100000001101100001111100110001010111111101111011011001011001001011100111101101111110100011011100100010001011111011001100000110011101010000100001001111101111011110000000100001101100100011100010101110001111010011010110110111011111110010100000111110011100011"
    );

  constant CIM_SEED : hypervector(0 to HV_DIMENSION-1) := (
		"1011111101111011110000100011001110100101101011100110100110001010011101110110001101001011110000000110000110010110010011001011000111110111100101110111101000000000000111000011010111111111001010100001110011101000010100111111111010011110111111011010100100110010000110010010110000000110011010001111011010000010001001010111100000001110111010110101101101000100110100011001110101110101101011001001101111101001010111101001000010101100001111000101001110100101001001101100011001101000001101110011111101111011011100010100101110001000010101011011101111101000001001110000100101001000110100000101000101110101001000001100101111010000100000000000111001000011101101000011000010101011101101001011010111101101101001111001011111101010011010000111011001111101101111101001100100001111000100001001001100101001111001111110110011100101001010000110011010111000001111100011111001000001000010001101000100101110000011010101011000000010110110101111101111010101110001011001001101000110110111001110000010110001111011100101101100100010010001001100100101000111"
    );

  constant IM_CONNECTIVITY_MATRIX : hypervector_array(0 to INPUT_CHANNELS-1)(0 to HV_DIMENSION-1) := (
		"1001101110010101000100000101101111110110111101011000110110100011101010100100100100001011000110110110010101100001111100000110111111100101000000000010111011011110111010001011010011100100001001010011101011010011010110011101000001011111000001001101110100101111110101000111010000010110101110100110111000110000000001110010001110010100100010100111111001011011000000000000000000000100101110011000110101110100000010100111001110011111001100100100000100101001100101010110101010110101011000110110000100111001110001111011010001101100000100011111110000000111001111111110110111010011011101110101110100000000010100010010000101111011110111000110101100011110000011101101010111001111101010111101101110010010010100100011001000001010010101010001000001111010111010100111010110100011000101010100000001101100001111100110001010111111101111011011001011001001011100111101101111110100011011100100010001011111011001100000110011101010000100001001111101111011110000000100001101100100011100010101110001111010011010110110111011111110010100000111110011100011",
		"0111001001110101101110001101001000000100100001010101100100110110001010111111111110011010101100100101110101010011000010001100100000011101100000000110100010010000100011011010011110011110011111011110001010011110010101110001100011010000100011111001000111101000000101101100011000110100101000111100100101101000000011001111011001110111110110111100000111010010100000000000000000001111101001110101100101000110000110111100111001110000111011111110001111101111011101010100101010100101010101100101001111100111001011000010011011001010001110110000001000001100111000000000100100011110010001000101000110000000110110111111001101000010000100101100101010110001000110001001010100111000001010100001001001111111110111110110111100011011110101011011100011000010100010111100010100110110101101010110000011001010011000011101011010100000001000010010111010111111010011100001001000000110110010011110111011010000010111010001101110001011001110011111000001000010001000001110011001011110110010110101001011000011110010100100100010000001110110001100001110010110",
		"1100111111000101001001011001111100001111110011010101011111100101011010100000000001110010101011111101000101011110100111011011110000110001010000001100110111111001110110010011110001110001110000010001011011110001110101001011010110011001110110000111101100001100001101001010110101100111101101100011111101001100000110111000010111000100000100100010001100011110110000000000000000011000001111000101011101101101001100100011100111001001100010000001011000001000010001010111101010111101010101011101111000011100111010100111110010111011011000101000011100011011100100000001111110110001111011101101101101000001100100100000111001100111001111101011101010101011101101011111010111100100011010110011111111000000000100000100100010110010000101010010010110100110110110100010110111100100101001010101000110111011110100110001010010110000011100111110100010100000011110010011111100001100101111110000100010011000110100011011001001011010111001110000100011100111011100011001110111010000101110100101111010100110001110111111110111000011000101011010011001110101",
		"0011100000101101111111010111000010011000001110010101010000011101010010110000000011001110101010000001101101010000111100010010001001101011011000011011100100000111000101111110001011001011001000111011010010001011000101111010010101110111000101001100001010011010011001111010100101011100001001010110000001111010001100100100110100101110001111110111011010110000101000000000000000110100011000101101010001001001111011110110011100111111010111000011010100011100111011010100001010100001010101010001000100110011100010111100001110100010010101101100110010110010011110000011000000101011000010001001001001100011011111110001100111011100111000001010001010101010001001010000010100011110110010101110000000100000001110001111110110101111001101011111110100111100100100110110100100011111101111010101101100100010000111101011011110101000110011100000110110110000110001111110000010011011101000001001110111110101100110110010111111010010100111001001110110011100010010110111000100011001101000111101000010111101011000100000000100100110101101010011110111000101"
    );

  constant CIM_CONNECTIVITY_MATRIX : hypervector_array(0 to INPUT_QUANTIZATION-2)(0 to HV_DIMENSION-1) := (
		"0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000100000000000100000000000000000000000100010000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000010001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000010000001000000",
		"0000000000000000000000000000001000001000000000000000000000000000000000000000000010000000000000000000000000000001000100000000000000000000000000000000000100010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100100000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000100000000011000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000",
		"0000000000000010000000000000000000000000000000010000000001000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010100000000000000010000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000100001000000000010000000000000000000000010000000000000000000000010000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000010000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000010010000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000011000000000000000100000000000000000000000000000000000000000000000000000000100000000010000000000010000000000000000000000000000000010001000000000100000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000010000010000000000000000000000000100000000000000000010000000000000000010000000000000000000000000000000000000000001000100000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000100000000000000000000000000010000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000110000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
		"0000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010001000000000100000000000000000000000100000000000000001000000000010000000100000010000000000000000000000",
		"0000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000100100000000100000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000101000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000001000000000000000000010000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"0001000000000000000000000000000000100000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000100000000000000000000000000000001000000000000000000010000000000100000000000000000000010000000000000000000000000000001000000000010010010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000010000000010000000000000000000100000000000000000000000000000000000000000000001000000000000110000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000",
		"0000000000000000000000000000000001000000100000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000010100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000010000000000000100001000000000001000000000000000000000000000000000000100000010100010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000",
		"0000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100100000000000000001000000000000000000000000001000000001010000000000000000000000000000000000000100000000000000000000000000000001000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000100000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"0100100000000000000000000000000000000000000000000000000000000000100000000000000000000001010000000000000000000000000000000000000000001000000000000000000000000000001000001010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000100000000001000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000001000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000100000000000100000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000001000000100000000000000000000000000000000000000000000000000000000000010000001010001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
		"0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000010000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000001000000001000010000000000000001000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000100000001000000001000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000010000000000001000000000000000000000000000000000001000000000000000000000000001000001000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000100000000000000000000000000000000010000000000000000010000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000001000001000000000000000000000000100000000000000000000000000000000000000000010000000000000000000010000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000",
		"0000000110000100000000000000000000000000000000000000000000000000010010000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000010000000010000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000100001000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000100000000000000000000000000100000000000000000000000000100000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000010000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001100000010000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000010000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
		"0000000000000000000000100000000000010000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000010000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000010100000000000000000000000000000010000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000001000000000000000000000000000000000000000101000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000010000000100000000000000000"
    );

  constant BUNDLE_CONNECTIVITY_MATRIX : hypervector_array(0 to MAX_BUNDLE_CYCLES-1)(0 to HV_DIMENSION-1) := (
		"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		"0001110111011100000111010000110100100110100111110001001010101110011001001010001010001001100101111010101100010011100101000001010101111001111000001100110100110000111000001111111010100110111010101011000001101010110001011001110010110010111100101101111100111010110100101010001000111010111001000011000110001000010111100100100110101011100101111101001011101011110101111100100100000011101100011010011111110001110000001101111101100001100100010000011110000001011010001111100010001010010100110011001010110011011000110100110111001111000101101000000110000011110111011110001110000110100100111101010011010100010000111100101110111100011001011010110000110110111000110010111100100110011011111010110010101101011001000011001110110010001011011001100010100100011011010111111001000000010010011100010101001110011100010101000001000110110100010001001111100111111001010101001111111011010101111100000100101111011011101000111101001101111110111011000010100110100010100110001110111000100000100111101110010111100110010110000001111011011100001101001010111011",
		"0001010000001000010110000001001000000001001010011000011000000000100000001100100010000101111000001100010100010001000011010001000000000100001001111110001100001001000101010000100011000011010010100111000001000001000100111101000010001000000110101100010100110000011010000001000001000100000000100010000010100010101100110000000111111100000101100000001100000100110000001001001110100110010000010000010001011010010111000010000011001000000000001011010000100011000000001000000000010001110000000001100000000001001101000011010010100100100100000010011000000000000100100000000000011000100000010000001100000010011110111101100001110110000000000011000011010000101100010011010110000111001000000000101000001011100000010010100000100011100100001010100000100000101001000000100011010110000000110000011100111000000001011001001111010010010011100000001111101000011001000010011101110101101100000101100010000010100010101001001010001000101011100100010011010111100011000000110000010010100000011100000100100000010000000011000101010000110110100100010000100010",
		"0010000110110000000000001111000000001110001000000001000100101000000001000000001000000011110001000110100101001000100101010100001000000000000100000000010010000000000000000111000000010000100000000001001001010001101010110000010011000101100000000001000000010010100000100000011001100001000000101000001010010101000000000000010001010000101100100000110010001000000110100000010000010010110100011100000000000101000100100000010011001010011000001110001001010010000110000000000000100000010111010000000001010000000001000000100000011100000101010010010001001001011000111010100000000000000000001000101001000000000100001000100011111000100000010000010001000000000100001000000010100110000000000110000000100100000000010001000001000110000100000001101000101010110100101010000100001000010000000000000010000001100010000100011000000000000000010001100000000010110011010100010100100111010000001000001010001011000000000000011100001100100001000110001000100001000110011000101000000000001010000010000100010000000000100100101000010110000010110011000000000000",
		"1110000000000010000001010000000000000000000000101000100000000010110100010011001000001100000000100100000100010000000000001001000000000000010000111000000010010000000000101000100000000000000000001000000001000100001100001001001000110000010010011010001100000001000000110001100000010011010000010000000000100011101100000100100100000010000010010100000100000001001011100000100100100000000000000000000000010000000110100000000010000100000000010001000001000000001000001001010000000011000100010000110100001100000000110000000000000010100000000000000010100000000100001001000000001000001110000000010000100000001001100000000000101100000000000011000001101010010001000100000011000000001000010000001000000000001011000010000000000101010001001000010100011000100001010000000000000010000001001101010100000000000001110000001000000011000000010011000001110000000100111100001000100000000100101100010000000010000000110000000000110000001000001100000010101000000000000000100001000000000000001000110010010101000000000000000000000100000001001000001000001101",
		"0000000000000000010001100000000000010000010010000000000100001101000001000001000000000101000000000010000100000000000100000000100000001010000000000000000100100111000000000000000010100000001000000000011000000000000000100001000000000110000011000010010000000010000001000100000001000000100001000000000010000000000010000001000010100010001000100000000010000001000000100000000100000001001100110001000010000010000000001000000010000000011001001000010000010100000000000000000000110000000001010100000000100100000000100000010000001000000000000000010000000010100010100001000011000010011000100000000000000000101000000100000010000100010100111000000100001000011000000001000000000100000000000000000000000000100000000010000010110001000110100000000001010010000000000001000001000101000101101010000100010000000000000001010000000000101000010010000000000000000000010000010001011010000100001010100000000000100100000001000010000101011010110000000100000010000110000000000000000101010100000100000000000000000000000000000010000000000011000000001000001000",
		"0010101000000000001000011000010000000000100000010001000000000000101000001000000000001000000010110100000000001010000000000010000000110101000100010000100011010010000011100000010100110000000000001000000000000100000011000100000000000000000110001000101000100000000000100000110000000010000000101000100000000000000010000000000101000010000000100101000110000010010000001000000000000111010000000100000100010000000000000000100000010000100100000001100000000000000000000000000000000010010000010000000000000000000000000000000010101000100000000110000000000100011000000100000000100000000000011100000110000000010011001100111010000000010000000001001000001000000000000000000100000000000000000000000010000010000000000010000011010000000000100000000000000000111000000000000100100100000000000000000010010000101000000000010000000000000000000100000100000000000001000000000010100001000001100000000000000001100001000010000010001000000100100000000100000001000000000100101000000101000000000001000000010000000000100100000000000101001000001000100000011000",
		"1000000000000001100010000000000001000000000010001000000000000010000000000000000000010000000011000000000000000101011000010011001000000010001001010000000000000000100000001010000000010000000000011000000000000000001000001000000000000000011000000000000000000000000000000000000000001000000001100101000000001000011000000001010001000000100000100000000000000000010000100000000010000001100000000100000000000000010010000000100000001101010010001000000000000000001000000000000000001010000010101100001101000000001001000000000100000010000000001000010000000000000010000001000000100000001010000000000000000000000101000000001100000001000000110001001010000000010001000010000000100000000100100010000001000101010000000000001000000000000000100010000001000000001000000000000000000000110000000000000000000000000000000001000000000000010110000000100000000000000001000000000000100000000000010000000000001000010000000000000010010000001010000000100000100010001010011000000001000001001011100000000000000000000000010001000000000100000000000000110000000000",
		"0000010000000100100000000000000000100110001000000000101000100001000000010000100000010100000000000000010000010000000000000000001000000000000000001000000000000011000000000001000000000001000001000000000001010000000000010000000010001000001000001001000010001000000100000000000100000100000000000000000000000000000000000001000000000000000000000001000010000000000000010000000100001000010000000000000000010000000000000000100000000000000010010000000000000000010000110000010000000000100000000000000000000000000010000000000101000000000100000000001100000010000000001010010000100010000101000000000000010000000000000000001000000000100000000000000001000000000000001000000000000000000010000100100000010010100000010000101100010010000100000000100000010000101000000000000000000000000000000000001000000000000000100000000001000000001001100000000000000101000010000000100000000000000000000101000010000000000000001000000000000000001010000000100010000010010000000000000000000000000010000000000000100000001000001000000000010110000000000100101000000000",
		"0000000000000010000010100000000000000000000000000000010000000000000001000000010011000100000001001000000000000100000001000000000001100100000000010001000000001000011000000000001000001000011110010000000100000000001000000000000100000000001100001000000010000000000000000100000000010000000000000000000000000100000000000100110010100110010000000000000000000000000000000001000000000000000000001000000000000000000000001000000000010000000000000000001000000000000001000000000000010001010010000000000100000000000000000000000100010000000000001101010000000001000000010100000000000000000000000000000000000000000000001000000000000001000001011000100000000011000100100000000010000100100000010000000000010000000000000100000000000000000000000000011000000000000000000000000000000000000001000000010100000000000000000000000000011100000000010000001000000001000000000000000000000000000000000000000000000000000000000000100000000010001010000010000000000000000010000000000100100001000000000001000100100000000000000001000010000000100100010001100000000100",
		"0000000000000000000000000000000100100000100000000000000001000000011000100000000000000000000000000101000000000001000000000000000000000100000000010000000000010000000000010000100010000000000000010000000000000000000010000101000000000000000000000000100000000000000000000000100000000000000100100000100000000100001000000000010000001000000000000000000000000100000000000001000010000000001000000000000000100001000000010100000000000000000000000100000010000000000000000000000000000000001000000000000100000010000000000100000010000000000000010000001000000000000001011010000011010001000000000100001000000001000000000000100000000000000100000000100101000010001000000010100100000010000000010000000000000000000100000000000000001000100000000000100000000000000000001001001000000000000000000000000000000000000000000000000000010000000000000010010000000000000000000000000000000100000000010000000001000000000100000000000001000010000000000000000000000000000000001000000000000001000000000000000010001000000000000000000000000100000000010000000000000010",
		"0010000000000000001011000010100010000100000000000001100000000000000000000000010010000000000000000000000000000000000010000010100000001000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000100000010000000000000000000000000100000100000100001000000000000000000000000000000000000001000000001000000000000000000000010000000000000001000010000000000000001000000001000000000000001000000000001000000000000001000000000000000000000000000100000010000000000000000000000000000000000000010000000000000100000000000000010000000110000001000000000000000000000000000001011000000000000000000000000000000000000000000010000010010000000000000000000001000001000000000000000000000001000000000000000000000000000000000000000000000000101011000000000010000000010011000010010000000000000000000000000100000000000010000010000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000100100000000000000010000000000000000000000100000000000000000000001010000000001001000000001000000000001000000000000000001000000000000010000000000000000010100000000010000000000010000000000000000000000000110000000000000001000000000000000100000000000000000000000000010000001010000000000000000100000010000000100000000000000001000001000000101000000000010000000000000000000000000000001000010000000010000000000000001000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000001000000000000000100000001100000000100001000000000000000000000001000000000000000101010000000000000000000000000000000000010000000000110000000000001010000000000000000001001000000000000000000000000000000000000000010011000000000000000000000000000011010000010000000000000000000100001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001000000001000001000000000001000000000000000000000000010000011000000010000000000000000000100010000000",
		"0001001000000000010000100000000000000000000001000000000000010000000000000000010000000000000000001100000010000000000000000000000000000000100000000101010000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000010000001000100100100100000000000000000000001000000010000000001000000000100000000010010000001001000000000000010000000000000010000010000000000000100010000000000000000000000000010001000000000000001000000000000000000010000001000000000000000000000000000011000000000000100000010001000000000000010000000000000010010000000000000001000000000000000000000000100000011100000000000000100000000000000010000000000000000000100000001000000000000000100000000000100000000000000010000000000000100000000010000000000000000000000011000000000000000000100000000100100000001000000000000000000000001000000100000010100000100000000000000000000000000100000000010000000000000000000000000000000001000010000000000001110000000000100001000010000000000000000000000000000000000000000000000000000000001",
		"0001000000000000100000000010000000000000000000000000000000000000001000000010001000000000000000000000000000000000000000010000000000010000000000100000100000000000000000000000000000000001000000000000000000000000000000000000000010000001000000000000000000000100000000100000100000011000000000000000000000000010010000000000010000010000000000000001000000010010000010000000000100010100000000000000000000001000000000000000000000000000000000000000000011000000000001000000000000000000001000000001000100000000000000010000000000000000000000000000100010000000000000100000000000000000001000000000000000100000000000001000001110000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000001010000000000000000000000000000000000000011000000000000001001000000000000000000000000000000001001100000000010000000000000000000000000000000000000000000000000000100000000000000000000001000000000101010000010000000010000001000000000000000000000",
		"0000000000000000010000000000000000000000010001000000000000000000000000000000000000100000000000000010000000000000000000000101000000000000000100000000000000000000000000000000010100000000000101000000000000010000000000000010000000001000010000000000000001000000000100000000000000000010000000000000000000000011001000000000000000001000000000000001100000000000010000110000000000000000000010000000010000010000000000000000000000000000000000100100000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000010000000000000000000110000000000000000000000000000000000100000000000000000000000000001000000000010001000000000000010000000000000010000000000000000000100000100000000100000000000000000000000001000000000000000000000000000001000000001100000000000010000000000000000000100000000000000",
		"0000000000100000100000000010000000000000000000000000100000010000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000001010000000000000001000000000000000000000001010000000000000000000000001000000000000000000000001000010000000000000000000000000000010001000000001010000000000000011000000000000000000000000000000000000000000000000000000110000000000000100000000000000000000000000000000000100000000000000010000000100001000000000011000000000010000000000000000000000000000000000000000000000000100000000000111000000100000100010000000000000000000100000000000000001000000000000010110000000000000000001000000000000100000000001100000010000000000000000000000000000000010000000000000000010000000000000000000000010000000000000000000000000000011000000000000000000000000000010001000001001000000000000000000000000000100000000000000010000000000100000010000100000010000000000000010100000000000100000000000000010100000000000000000000000000000000000000000000000100000000",
		"0000000010100001001000000000001000000000000000000000000000010000100000100000000001000100000000000000010000000000000000000010000000001000000001001100000000000000000000000000000000000000000010000000000000000000100000000000001010000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000001000000000000000000100110000001000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000010000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000100000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001001000010001000000000000000000000001000000000010000000000100000000000000000000000000000001000000000001000000000000001000000001000000000000000001000000000001000000000100000000100000000000010100000100000000000010000000000000000000000000100000001000000000010000000000000000000000000",
		"0000000000001000000000000100000000000000000000000000000110001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000100000000000000000100100000000000000000000000000000000000000100000100000000000000000001001000000000000000000010000000000000100000000000010000000000000010000000000001000000000000000000000100001110000100000100000000000000000000100000000000001000000000000000000000001010000000000000000001000000000000000000000000010000000000000000000000001000000001000000000000000000000000100000000000000000000000000000000000000010000000000000000001000000000000000000100000000000010000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000100000000000001000001000000000000000000000000000000000000000000000000000010000000000000000010100000000000000000000000000000001000000000000000110000100000011000000000000000000000000000000000000000000000000000001000000000000110000000000001000000000010000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000001000000000000000000010100000000100000000000000010000000000000000000000100000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000001000000000000000001010000000000000000000000000000000000000000000000000100000000000000001100000000000001000000000100000000000000000000001000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000010010000000000000100000001000000000000000000100000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100000000000010000000000000000000000000000001000000010100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000",
		"0000000000000000000001100000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000010000000000000000100000001000000000001001000000000000000010000000000000000000000000100010000100100000000000000000000000000000000000001000000000000000000001000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000100000001000100000000000100100000000001000000000100000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000100000000000000000000100000000100000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000100000001000000000000000000000001001000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100000000011000100000000000000000000000001000000000000000010000000000000000000000010000000000000000000000000001000000000000000000000000",
		"0000000010000000000000000010000000100000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000100000000010000000100000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000001000000000101000000100000000100010000000000000000001000000000000000000000000000000000000000000001000100000000101000100000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000101100000000000000100000000000000000000000000000000000000000000100000000001000000010000000000000000000000000010000000000000000000000000000000000100000000110111000000000100000000000",
		"0000000001000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000001000000000000100000000000000000000000000100000001000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000100000000001100000000100010000000000100000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000001000000000000100000000000000100000000000000000000000000000000000000000000100000000000000010000000100000000000000000000000000000001000000000000000000000000000000000000000000000000010000100000000000100000000",
		"0000000000000000010000000100001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000110000000000010000000000000000000000000000000000000000100000000000000000000010000000000010000000000000000000000000000000011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000010000000000000000010010100000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000010000000000000000000000000000000000000000000100000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000010000000000",
		"0000000000100001000000000010000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000001000000000000000010000001000000000000000000000100001000000000000000000001000100000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000010000100000000000000000000010000000000000000000010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000100000000000000000000000000000001001000000000000000000100000000000000000000010000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000",
		"0000000000000000001000000000000001000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000010010000001000000000000000000000000000000000000010000000110000000000101000000000000000000000000000000001000000000000000000000000010010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000100000000011000000000000000000001000000000000000000000000100000000000000000000000100100000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
		"1000000000000100000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010010000001000000000000000000100000001000000000000000010001000000000001000000000000000000100000000000000000000000000000000000000000101000001000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100010000000000000000000000000000000000100001000000000000000000000000000000000000000000001000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000100000000000000100000000000000000000000000000000000000000100000000000000000000000000000000001101000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000010000000001000000000000000000000000000000000000000000000000100000000000000000001000000100000000000000001000100000000000000000000010000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000001000000001000000000001000000000000000000000000000000000000100000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000100000000000000000000000000000001000000000000000000000",
		"0010000000000001000000000000001000000000000000010000000000000000001010000000000000000000000000000100000100000000000000010000000000000000000000000000000000100000000000000000000001001000000000000000000000000000000000000000100000001000000001001000000000010000000000000110000000000000000000000000000000000000000000001000000000010000000000000000000000000001000000000000000000000001001000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000010000000000000000100000000001000000001000000000000000000000000010000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000",
		"1000000001000000000000000100100000000000000000010000000000000000000010000000000000000000000000000000000000100000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000110000000000010000000010000000000000000000000000000000000000000000100010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000100000100000000000000010000000000000000000010000000000000000000000000100000000000000010000000000000000000000000000000000000010000000000100000001001000000000000000000000000000000000100000000000000000000000000000000010000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000001010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000010000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000100000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000",
		"1000000000000000000000000000010000000000001000000000000010000000000000000001000000100000001000000000000001010000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000001000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000100000001000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000100000000000000010000000000"
    );

end hdc_enhanced_pkg;

-------------------------------------------------------------------------------

package body hdc_enhanced_pkg is

  

end hdc_enhanced_pkg;

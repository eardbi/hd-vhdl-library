-- Copyright 2018 ETH Zurich
-- Copyright and related rights are licensed under the Solderpad Hardware
-- License, Version 0.51 (the “License”); you may not use this file except in
-- compliance with the License.  You may obtain a copy of the License at
-- http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
-- or agreed to in writing, software, hardware and materials distributed under
-- this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
-- CONDITIONS OF ANY KIND, either express or implied. See the License for the
-- specific language governing permissions and limitations under the License.

------------------------------------------------------------------------------
-- Title      : HDC Baseline Package
-- Project    : Semester Thesis I
-------------------------------------------------------------------------------
-- File       : hdc_baseline_pkg.vhd
-- Author     : Manuel Schmuck <schmucma@student.ethz.ch>
-- Company    : Integrated Systems Laboratory, ETH Zurich
-- Created    : 2017-09-30
-- Last update: 2018-01-02
-- Platform   : ModelSim (simulation), Vivado (synthesis)
-------------------------------------------------------------------------------
-- Description: Provides the memories and functions required by the
--              baseline architecture.
-------------------------------------------------------------------------------
-- Copyright (c) 2017 Integrated Systems Laboratory, ETH Zurich
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author    Description
-- 2018        1.0      schmucma  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.hdc_pkg.all;

-------------------------------------------------------------------------------

package hdc_baseline_pkg is

  -----------------------------------------------------------------------------
  -- Function Declarations
  -----------------------------------------------------------------------------
  function majority (hvarray : hypervector_array) return hypervector;

  -----------------------------------------------------------------------------
  -- Constant Declarations
  -----------------------------------------------------------------------------
  constant ITEM_MEMORY : hypervector_array(0 to INPUT_CHANNELS-1)(0 to HV_DIMENSION-1) := (
		"1001101110010101000100000101101111110110111101011000110110100011101010100100100100001011000110110110010101100001111100000110111111100101000000000010111011011110111010001011010011100100001001010011101011010011010110011101000001011111000001001101110100101111110101000111010000010110101110100110111000110000000001110010001110010100100010100111111001011011000000000000000000000100101110011000110101110100000010100111001110011111001100100100000100101001100101010110101010110101011000110110000100111001110001111011010001101100000100011111110000000111001111111110110111010011011101110101110100000000010100010010000101111011110111000110101100011110000011101101010111001111101010111101101110010010010100100011001000001010010101010001000001111010111010100111010110100011000101010100000001101100001111100110001010111111101111011011001011001001011100111101101111110100011011100100010001011111011001100000110011101010000100001001111101111011110000000100001101100100011100010101110001111010011010110110111011111110010100000111110011100011",
		"0111001001110101101110001101001000000100100001010101100100110110001010111111111110011010101100100101110101010011000010001100100000011101100000000110100010010000100011011010011110011110011111011110001010011110010101110001100011010000100011111001000111101000000101101100011000110100101000111100100101101000000011001111011001110111110110111100000111010010100000000000000000001111101001110101100101000110000110111100111001110000111011111110001111101111011101010100101010100101010101100101001111100111001011000010011011001010001110110000001000001100111000000000100100011110010001000101000110000000110110111111001101000010000100101100101010110001000110001001010100111000001010100001001001111111110111110110111100011011110101011011100011000010100010111100010100110110101101010110000011001010011000011101011010100000001000010010111010111111010011100001001000000110110010011110111011010000010111010001101110001011001110011111000001000010001000001110011001011110110010110101001011000011110010100100100010000001110110001100001110010110",
		"1100111111000101001001011001111100001111110011010101011111100101011010100000000001110010101011111101000101011110100111011011110000110001010000001100110111111001110110010011110001110001110000010001011011110001110101001011010110011001110110000111101100001100001101001010110101100111101101100011111101001100000110111000010111000100000100100010001100011110110000000000000000011000001111000101011101101101001100100011100111001001100010000001011000001000010001010111101010111101010101011101111000011100111010100111110010111011011000101000011100011011100100000001111110110001111011101101101101000001100100100000111001100111001111101011101010101011101101011111010111100100011010110011111111000000000100000100100010110010000101010010010110100110110110100010110111100100101001010101000110111011110100110001010010110000011100111110100010100000011110010011111100001100101111110000100010011000110100011011001001011010111001110000100011100111011100011001110111010000101110100101111010100110001110111111110111000011000101011010011001110101",
		"0011100000101101111111010111000010011000001110010101010000011101010010110000000011001110101010000001101101010000111100010010001001101011011000011011100100000111000101111110001011001011001000111011010010001011000101111010010101110111000101001100001010011010011001111010100101011100001001010110000001111010001100100100110100101110001111110111011010110000101000000000000000110100011000101101010001001001111011110110011100111111010111000011010100011100111011010100001010100001010101010001000100110011100010111100001110100010010101101100110010110010011110000011000000101011000010001001001001100011011111110001100111011100111000001010001010101010001001010000010100011110110010101110000000100000001110001111110110101111001101011111110100111100100100110110100100011111101111010101101100100010000111101011011110101000110011100000110110110000110001111110000010011011101000001001110111110101100110110010111111010010100111001001110110011100010010110111000100011001101000111101000010111101011000100000000100100110101101010011110111000101"
    );

  constant CONTINUOUS_ITEM_MEMORY : hypervector_array(0 to INPUT_QUANTIZATION-1)(0 to HV_DIMENSION-1) := (
		"1011111101111011110000100011001110100101101011100110100110001010011101110110001101001011110000000110000110010110010011001011000111110111100101110111101000000000000111000011010111111111001010100001110011101000010100111111111010011110111111011010100100110010000110010010110000000110011010001111011010000010001001010111100000001110111010110101101101000100110100011001110101110101101011001001101111101001010111101001000010101100001111000101001110100101001001101100011001101000001101110011111101111011011100010100101110001000010101011011101111101000001001110000100101001000110100000101000101110101001000001100101111010000100000000000111001000011101101000011000010101011101101001011010111101101101001111001011111101010011010000111011001111101101111101001100100001111000100001001001100101001111001111110110011100101001010000110011010111000001111100011111001000001000010001101000100101110000011010101011000000010110110101111101111010101110001011001001101000110110111001110000010110001111011100101101100100010010001001100100101000111",
		"1011111101111011110000100011001110100101101011100110100110001000011101110110001101001011110000000110000010010110010011001011000111110111100101110111101000000000000111000011010111111111001010100001110011101000010100111011111010011110111110011010100100110010000110010010110000000110011010101111011010100010001001010111100000101100111010110101100101000100110100011001110101110101101011001001101111101001010111101000000010101100001111000101001110100101001011101100011001101000001101110011111101111001011100010100101110001000010100011011101111101100001001110000100101001000110100000101000101110101001000001100101111010000100000000000101001000011101101000011000010101011101101001011010111101100101001111001011111101010011010100111011001111001101111101001100100001111000100001001001100101001111001111110110011000101001010000110011010111000001111100011111001010001000010001101000100101100001011010101011000000010110110101111101111010100110001011001001101000110110111001110000010110001111011100101101000100010010001001110100100000111",
		"1011111101111011110000100011000110101101101011100110100110001000011101110110001111001011110000000110000010010111010111001011000111110111100101110111101100010000000111000011010111011111001010100001110011101000010100111011111010011110111110011010100100110011000110010010110000000110011010101111011010100010001001010011000000101100111010110101000101000100110100011001010101110101101011001001101111101001010111101000000010101100001111000101001110100001001011101100011001101000001101110011111101111001011100010100111110001000010100011011101111101100001001110000100101001000110100001101000101110101000000001100101111010000100000000000101001000011101101000011000010101011101101001011010111101100101001111001011111101010011010100111011001111001101111101001100100001111000100001001001100101001111011111110110011000100001010000110011010111000001111100011111001010001000010001001000100110100001011010101011000000010110110101111101111110100110001011001001101000110110111001110000010110001111011100101101000100010111001001110100100000111",
		"1011111101111001110000100011000110101101101011110110100111001000011101110110001111011011110000000110000010010111010111001011000011110111100101110111101100010000000111000011010011011111001010100001110011101000010100111011111010011110111110011011100100110011000110010010110000000110011010101111011010100010001001010011000001100100111010110101000101000100110100011001010101110101101011001001101111101001010111101000000010101100001011000101001110100001001011101110111001101000001111110011111101111001011100010100111110000000010000011011101111101100001001110000100101001000110100001101000111110101000000001100101111010000100000000100101001000011001101000011000010101011101101001011010111101000101001111001011111100010011010100111011001111001101111101001100100001111000100001001001100101001111111111110110011010100001010000110011010111000001111100011111001010001000010001001000100010100001011010101011000000010110110101111101111110110110001011001001101000110110111001110000010010001111011100101101000101010111001001110100100000111",
		"1011111101111001110000100011000110101101101011110110100111001000011101110110001111011111110000000010000010010111010111001011000011110111100101110111101100010000000111000011011011011111001010100001110011101000010100111011111010011111111110011011000101110011000100010010110000000110011000101111011010100010001011010011000001100100011010110101000101001100110100011001010101110101101011001001101111101001010111101000000010101100001011000101001110100001001011101110111001101000001111110011111101111001011100010110111110000000010000011011101111111100001001110000110101001000110110001111000111110101000000001100101111010000100000000100101001000011001101000011000010101011101101000011010111101000101001111001011111100010011010100111011001111001101111001001100100011101000100001001001101101001111111111110110011010100001010000110011010111000001101100011111001011001001010001001000100010100001011010101011000000010110110101111101111110110110001011001001101000110110111001110000010010001111011100101100000101010111001001110100100000111",
		"1011111101111001110000100011000110101101101011110110100111001000011101110110001111011111110000000010000010010111010111001010000011110111100111110111101100010001000111000011011011011111001010100001110011101000010100111011111010011101111110011011000101110011000100010010110000000110011000101111000010100010001011110011000001100100011010110101000101001100110100011001010001110101111011001001111111101001010111101000000010101110000011000101101110100001001011101110111001101101011111110011111101111001011100010110111110000000010000011011101101111100001001110000110101001000110110001111000111110101000001000100101111011000100000000100101001000011001101000011000010101011101101000011010111101000101001111001011111110010001010100111011001111001101111001001100100011101000100001001001101101001101111111110110011010100001010000110011010111000001101100011111001011001001010001001000100010100001011010101011001000010111110101111101111100110110001011001001101000110110111001110000010010001111011100101100000101010111001001110100100000111",
		"1011111101111001110000110011010110101101101011110110100011001000011101110100001111011111110010000010000010010111010111001010000011110110100011110111101100010001000111000011011011011011001000100101110011101000010100111011111010011101111110011011000101110011000100010010110000000110011000101111000010100010001011110011000001100100011010110101010101001100110000011001010001110101111011001001111011101001010111101000000010111110000001000101101110100001001011101110111001101101011111111011111101111001011100010110111110000000010000011011101101111100001001110000110101001000110110001111000111110101000001000100101111011000100000001100101001010011001101000011000010101011101011000011010111101000101001111001111111110010001010100111011001111001101111001001100100011101000100001001001101101001101111111110110011010110001010000110011010111000001101100011111001011001001010001001010100010100001011010101011001000010111110101101101011100110110001011001001101000110110111001110000010010001111011100101100000101010111001001110100100001111",
		"1011111101111001110001110011010110101111101011110110100011001000011101110100001111011111110010000010100010010111010111000010000001110110100011110111101100010001000111000011011011011011001000100101100011101000010100111011111010011101111110011011000101110011000100010010110010000110011000101111000010100010001011110011000001100100011010110101010101001100110000011001010001110101111011001011111011101001010111101000000010111110000001000101101110100001011011101110111001101101011111111011111101011001011100010110111110000000110000011011101101111100001001110000110101001000110110001110000111110101000001000100101111011000100000001100101001010011001101000011000010101011101011000011010111101000101001111001111111110010001010100111111001111001101101001001100100011101000100001001001101101001101111111110110011010110001010000110011010111101001101100011111001011001001010001001010100010100101011010101011001000010111110101101101001101110110001111001001101000110110111101110000010010000111011100111100000001010101001001110100100001111",
		"1011111101111001110001110001010110101111100011110110100011001000011101110100001111011111110010000010100010010111010111000010000001110110100011110111111100010001000111000011011011011011001000100101100011101000010100111011111010011101111110011011000101110011000100010010110010000110011000101111000011100010001011111011000001100100011010110101010101001000010000011101010001110101111011001011111010101001010111101000010010111110000001000101101110100001011011101110111011101101011111111011111101011001011110010011111110000000110000011011001101111100001001110000110101001000110110001110001111110101000001000100101111011000100000001100101001010011001101000010000010101011101011000011010111101000101001111001101111110011001010100111111001101001101001011001100100011101000100001001001101101001101111111110110011010110001010000110011010111101001101100011111001011000001010001001010100010100101011010101010001000010111110101101100001101010110001111001001101000110110111101110000010010000111011100111100000001010101001001110100100001111",
		"1010111101111001110001110001010110001111100011110110100011000000011101111100001111011111110010000010100010010111010111000010000000110110110011010111111100010001000111000011011001011011001000100101100011101000010100111011111010011101111100011011000101110011000100010010110010000110011000101111000011100010001011111011000001100100011010110101010101001000010000011101011001110101111011001011111010101001010111101000010010111110000001000101101110101001011011101110111011101101011111111011111101011001011110010011111110000000110000011011000101111100001001110000110101001000110110001110011111110001000001000100101111011000100001001100101001010011011101000010100010101011101011000001010111101000101001111001101110110011001000110101111001101001101001011001100100011101000100001001001101101001101111111110111011010110001010001110011010111101001101100011111001011000001010001001010100010100101011010101010001000010111110101101100001101010110001111001001101000110110011101110000010010000111011100111100000001010101001001110100100001111",
		"1010111101111001110001110001010110001111100011110110100011000000011101111100001111011111110010000010100010010101011111000010000000110110110010010111111100010001000111000011011001011011001000100101100011101000010100111011101000011101111100011011000101110011000100010010110010000110011000101111000011100010001011111011000001100100011010110101010101001000010000011101011001110101111011101011111010101011010111101000010010111110000001000101101010101001011010101110111011101101011111111011111111011001011110010011111110000000110000011011000101011100001001110000110101001000110110001110011111111001000001000100101111011010100001001100101001010011010101000010100010101011101011000001010111101000101001111001101110110011001000110101111001101001100001011001000100011101000100011001001111101001101111111110011011010110001010001110011010111101001101100010111001011000111010101001010100010100101011000101010001000010111110101101100001101010110001111001001101000110110011101110000010010000111011100111100000011010101001011110100100001111",
		"1010111101111001110001110001010111001111000011010110100011000000011101111100001111011111110010000010100010010101011101000010000000110110110010010111111100010001000110000011011001011011001000100101100011101000010100111011101000111101111100011011000101010011000100010010110010000110011000101111000111100010001011111011000001100100011010100001010101001000010000011111011001110101111011101011111010101011010111101000010010111110000001000101101010101001010010101110111011101101011111111011111111001001011110010011111110000000110000011011000101011100001001110000110101001000110110001110011111111001000001000100101111011010100001001100101001010011010101000010100010101011101011000001010111101000101001111001101110110011001000110101111001101001100001011001000100011101000100011001001111111000101111101110011011010010000010001110010010111101001101100010111001011000111110101011110110010100101011000101010001010010111110101101100001101010110001111001001101000110110011101110000010010000111011100111100001011010101001011110100100011111",
		"1010111101111001100101110001010111001111000011010110100011000000011101111100001111011111110010000010100010010101011101000010000000110110110010010111111100010001000110000011011001011011001000100101100011101000011100111011101000111101111100011011000101011011000100010010110010000110011000101111000111100010001011111011000001100101011011100001010101001000010000001111011001110101111011101011111010101011010111101000010010111110000001000101101011101001010010101110111111001101011111111010111111001001011110010011110110000001100000011011000101011100001001110000110001001000110110001110011111111000000011000100101111011011100001001100101001010011010101000010100010101011101011000001010111101000101001111001100110110011001000110101111001101001100000011001000100011101000100011101001111111000101111001110011011010010000010001010010010111101001101100010111001011000111110101011110110010100101010000101000001010010111110101101100001101010110001111001001101000110110011101110000010010000111011100111100001011010101001011110100100011111",
		"1110011101111001100101110001010111001111000011010110100011000000111101111100001111011110100010000010100010010101011101000010000000111110110010010111111100010001001110001001011001011011001000100101100011101000011100111011101000111101111000011011000101011011000100010010110010000110011000101111000111100010001011111011000001100101011001100001010101001000010000001111011001110101111011101011111010111011010111101000010010111110000001000101101011001001010010101110111111001101011111111010111111001001011110010011110110000001100000011011000101011100001001110000110001011000110110001110011111101000000011000100101111011011100001001100101101010011010101000010100110101011100011000001010111101000101001111001100110110011101000110101110001101001100000011001000100011101001100011101001111111000101111001110011011010010000010001010010010001101001101100010111001011000111110101011110110010100101010000101000001010010111110101101100001101010111001111001001101000110100011101010000010010000111011100111100001011010101001011110100100011111",
		"1110011101111001100101110001010011001111000011010110100011000000111101111100001111011110101010001010101010010101011101000000000000111110110010010111111100010001001110001001011001011011001000100101100011101000011100111011101000111101111000011011000101011011000100010010110010000110011000101111000111100010001011111011000001100101011001100001010101001000010000001111011011110101111011100011111010111010010111101000010010111110010001000101101011001001010010101110111111001101011111111010111111001001011110010011110110000001100000011011000001011100001001110000110001011000110110001110011111001010000011000100101111011011100001001100101101010011010101000110100110101111100011000001110111101000101001111001100110110011101000110101110001100001100000011001000100011101001100011101001111111000101110001110011011010010010010001010010010000101001001100010111001011000111110101011110110010100101010000101000011010011101111101101100001101010111001111001001101000110100011101010000010010000111001100111100001011010101001011110100100011111",
		"1110010101111001100101110001010011001111000011010110100011000000111101111100001111011110101010001010101010010101011101000000010000111110110010010111111100010011001110001001001001011011001000100101100011100000011100111011001000111101111000011011000101011011000100010010110010000110011000101111000111100010001011101011000001100101011001100001010101001000010000001111011011100101111010100011111010111010110111101000010010111110010001000101101011001001010010101110111111001101011111111010111111001001011110010011110110000001100000011011000001011100001001100001110001011000110110001010011111001010000011000100101111111011100001001100101101010011010101001110100111101101100011000001111111101000101001111001100110110011101000110000110001100001100000011001000100011101001100011101001111111000101110001110011011010010010010001010010110000101001001100010111001011000111110101011110110010100101110000101000011010011101111101101100001101010111101111001001101000010100010101010001010010000111001100111100001011010101001011110100100011111",
		"1110010101111001100101110001010011001111000011010110100011000000111101111100001111011110101010001010101010010101011101000000010000111110110010010111111100010011001110001001001001011011001000100101100011100000011100111011001000111101111000011111000101011011000101010010100010000110010000101111000111100010001011101011001001100101011001100001010100001001010000001111011011100101111000100011111010111010110111101000010010111110110001000101101011001001010010101110111111001101011111111010111111001001011110010011110110000001100000011111000001011100001001100001110011011000010110001010011111001010000011000110101111111011100011001100100101010011010101001110100111101101100011000001111111001000101001111001100110110011101000110000110011100001100000010001001100011101001100011101001011111000101110001110011011010010010010001000010110000101001001110010101001011000111110101010110110010100101110000101000011010011101111101101100001101010111101111001000101000010100010101010001010010000111001100111100001011110101001011110100100011111",
		"1110010011111101100101110001010011001111000011010110100011000000101111111100001111011100101010001010101010010101011101000000010000011110110010010111111100010011001110001000001001011001001000110101100011100000001100111011001000101101111000011111000101011011000101010010100010000110010000101111000111100010001011101011001001100101011001101001010100001001010000001111011011100101110000100011111010111010110111101000010010111110110001000100101011001001010010101110111111001101011011111110110111001001011111010011110110000001100000011111000001011100001001100001110011010000010110001010011111001010000011000110101111111011100011001100100101010011010101001100100111111101100011000001111111001000101001111001100110110011101000110000110011100001100000010001001100011101001100011101001011111000101110001110011011010010010010001000110110000101001000110010101001011000111110101010110110010100101110000101000011010011101111101101100001101010111101111001000101000010100010101010001000010000111001100111100001011110101001011110100100011111",
		"1110010011111101100101110001010011001111000011010110101011000000101011111100001111011100101010001000101010010101011101000000010000011110110010010111111100110011001110001000001001011001001000110101100011110000001000111011001000101101111000111111000101011011000101010110100010000110010000101111000111100011001011101011011001100101011001101001010100001001010000001111011011100101110000100011111010111010111111101000010010111010110001000100111011001001010010101110101111001101011011111110110111001001011111010011110100000001100000011111000001011100001001100001110010110000000110001010011111001010000011000110101111111011100011001100100101010001010101011100100111111101100011000001111111011000011001111001100110110011101000110000110011100001100000010001001100011101001100011101001011111000101110001110011011010010010010001000110110000101001000110010101001011000111110101010110110010100101110000101000011110011101111101101100001101010111101111101000101000010100010101010001000010000111001100011100001011110101001011110100100011111",
		"1110010011111101100101010001010011011111000011010110101011100000101011111100001111111100101010001000101010010101011101000000010000011110110010010101111100110011001110001000001001011001101000110101100010110000001000111011001000101101011000111111000101011011000101010110100010000110010000101111000101100011001011101011011001100101011001101001010100001001010000001111011011100101110000100011111010111010111111101000010010111010110001000100111011001001010010101110101111001101011011111110110111001001011111010011010100000001100000111111000001011101001001100001110010110000000110001010011111001010000011000110001111111011100011001100100101110001010111011100100111111101000011000001111111011000011001111001100110110011101000110000110011100001100000010001001100011101011100011101001011111000101110000110011011010010010010001000110100000111001000110010101001011000111110100010110110010100101110000101000011110011101111101101100001101010011101111101010001000010100010101010001000010010111001100011100001011110101001011110100100011111",
		"1110010011111101100101010001010011011111000011010100101001100000101011111100001111111100101010001000101010010101011101000100010000011110110010010101111100110011001110001000001001010001101000010101101010110000001000111011001000101101011000111111000101011011000101010110100010000110010000101111000101100011101011101011011001100101011001101001010100001001011000001111011011100111110000100011111010111010111111101000010010111010110001001100111011001001010010101110101111001101011011111110110111001001011111011011010100000001100000111111000001011111101001100101110010110000000110001010011111001010000011000110001111111011100011001100100101110001010111011100100111111101000011000000111111011000011001111001100110010011101001110000110011100001100000010001001100011000011100011111001011111000101110000111011011010010010010001000110100000111001000110010101001011000111110100010110111010100101110000101000011110011101111101101100001101010011101111101010001010010100010101010001000010010111001100011110001011100101001111110100100011111"
    );

end hdc_baseline_pkg;

-------------------------------------------------------------------------------

package body hdc_baseline_pkg is

  -----------------------------------------------------------------------------
  -- Function Definitions
  -----------------------------------------------------------------------------

  function majority (hvarray : hypervector_array) return hypervector is
    variable sum    : integer                          := 0;
    variable result : hypervector(0 to HV_DIMENSION-1) := (others => '0');
  begin
    sum := 0;
    for i in 0 to HV_DIMENSION-1 loop
      sum := logic_to_integer(hvarray(0)(i));
      for j in 1 to hvarray'high loop
        if hvarray(j)(i) = '1' then
          sum := sum + 1;
        else
          sum := sum - 1;
        end if;
      end loop;  -- j
      if sum > 0 then
        result(i) := '1';
      else
        result(i) := '0';
      end if;
    end loop;  -- i
    return result;
  end majority;

end hdc_baseline_pkg;
